#define DES_ECB_DES_ECB_STR_ADDR 0
#define DES_ECB_DES_ECB_END_ADDR 0
#define DES_ECB_DES_ECB_CACHE_NUM 4

rcm_mem_rlm_array='{
0xc0200400 0x00000000 0x00000000 0xffff4000
};

rcm_mem_rcu_array='{
32'h00000000,32'h00048008,32'h00041800,32'h00000000,32'h00000000,32'h00000000,32'h0000fe00,32'h00000000,
32'h00000041,32'h02038008,32'h00031000,32'h00000000,32'h00000000,32'h00000000,32'h0000fe03,32'h00000000,
32'h00000042,32'h01028008,32'h41020800,32'h00030000,32'h02800000,32'h80401808,32'h0000fe00,32'h00000000,
32'h00200000,32'h00000000,32'h00008000,32'h00000000,32'h00000000,32'h00000000,32'h0000fe00,32'h00000000
};

rcm_mem_bfu_array='{
32'he0000010,32'h0003ffff,32'h00000000,32'h00000000,
32'h00000028,32'h0003fa8c,32'h00000000,32'h00000000,
32'h20000028,32'h0003fa9c,32'h00000000,32'h00000000,
32'h10906004,32'h0003f820,32'h00000000,32'h00000000,
32'h10014004,32'h0003f942,32'h00000000,32'h00000000,
32'h0000002a,32'h000162d4,32'h00000000,32'h00000000,
32'h80000009,32'h0003fad5,32'h00000000,32'h00000000
};

rcm_mem_route_array='{
32'h0fffffff,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd62d,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd021,32'h00000000,32'h00000000,32'h00000000,
32'h0fffc284,32'h00000000,32'h00000000,32'h00000000,
32'h0fffff86,32'h00000000,32'h00000000,32'h00000000,
32'h0fffc488,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd62c,32'h00000000,32'h00000000,32'h00000000,
32'h0fffc080,32'h00000000,32'h00000000,32'h00000000,
32'h0fffdebc,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd0a0,32'h00000000,32'h00000000,32'h00000000
};

rcm_mem_mem_ctrl_array='{
32'h00000001,32'h00000000,32'h000001e0,32'h00000020,
32'h00000001,32'h00000000,32'h200001e0,32'h00000000,
32'h00000001,32'h00000000,32'h020001e0,32'h00000020
};

