
`define twofish_STR_ADDR 0
`define twofish_END_ADDR 0
`define twofish_CACHE_NUM 4
rcm_mem_array='{
32'hc0200400,32'h00000000,32'h00000000,32'hffff4000
};
rcm_mem_rcu_array='{
32'h00000000,32'h00009908,32'h00000000,32'h08000000,32'h02008020,32'h82c0b830,32'h0000000a,32'h00000000,
32'h00000041,32'h02000000,32'h04000000,32'h28030001,32'h08824098,32'h81c07820,32'h00000006,32'h00000000,
32'h00000002,32'h01011908,32'h00000000,32'h18000000,32'h04814058,32'h80c03810,32'h00000002,32'h00000000,
32'h00100000,32'h00000000,32'h00000000,32'h08000000,32'h02008020,32'h00201006,32'h00000000,32'h00000000
};

rcm_mem_bfu_array='{
32'h00000028,32'h0003fae5,32'h00000000,32'h00000000,
32'h20000028,32'h0003faf5,32'h00000000,32'h00000000,
32'h40000028,32'h0003fac5,32'h00000000,32'h00000000,
32'h60000028,32'h0003fad5,32'h00000000,32'h00000000,
32'he0000010,32'h0003ffff,32'h00000000,32'h00000000,
32'h00000010,32'h0003fa89,32'h00000000,32'h00000000,
32'h00000010,32'h0003fa99,32'h00000000,32'h00000000,
32'h51010404,32'h0003fff9,32'h00000000,32'h00000000,
32'h00000010,32'h0003f850,32'h00000000,32'h00000000,
32'h40000010,32'h0003f840,32'h00000000,32'h00000000,
32'hd101fc24,32'h000267f0,32'h00000000,32'h00000000,
32'h10c20004,32'h0003fcd1,32'h00000000,32'h00000000,
32'hc0000009,32'h0003fcf9,32'h00000000,32'h00000000,
32'h00000028,32'h0003f912,32'h00000000,32'h00000000,
32'h40000028,32'h0003f932,32'h00000000,32'h00000000,
32'h80000028,32'h0003f952,32'h00000000,32'h00000000,
32'hc0000028,32'h0003f972,32'h00000000,32'h00000000,
32'h00000028,32'h0003f820,32'h00000000,32'h00000000,
32'h80000028,32'h0003f860,32'h00000000,32'h00000000,
32'hc0000009,32'h0003faf5,32'h00000000,32'h00000000,
32'h80000009,32'h0003fad5,32'h00000000,32'h00000000,
32'h80000028,32'h0003fa87,32'h00000000,32'h00000000,
32'ha0000028,32'h0003fa97,32'h00000000,32'h00000000,
32'hc0000028,32'h0003faa7,32'h00000000,32'h00000000,
32'he0000028,32'h0003fab7,32'h00000000,32'h00000000
};

rcm_mem_route_array='{
32'h0fffffff,32'h00000000,32'h00000000,32'h00000000,
32'h00c10100,32'h00000000,32'h00000000,32'h00000000,
32'h01e3860a,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd6ac,32'h00000000,32'h00000000,32'h00000000
};

rcm_mem_mem_ctrl_array='{
32'h00000001,32'h00000000,32'h1e0001e0,32'h00000000,
32'h00000001,32'h00000000,32'hfe0001e0,32'h00000001,
32'h00000001,32'h00000000,32'hfe0001e0,32'h00000007
};
