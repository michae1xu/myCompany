
`define TWO_FISH_STR_ADDR 0
`define TWO_FISH_END_ADDR 0
`define TWO_FISH_CACHE_NUM 4
rlm_mem_array='{
32'hc0200400,32'h00000000,32'h00000000,32'hffff4000
};
rcm_mem_rcu_array='{
32'h00000000,32'h00009908,32'h00000000,32'h08000000,32'h02008020,32'h00201006,32'h00000000,32'h00000000,
32'h00000041,32'h01000000,32'h04000000,32'h18020001,32'h04814058,32'h80c03810,32'h00000002,32'h00000000,
32'h00000002,32'h02019908,32'h00000000,32'h08000000,32'h08824020,32'h81c07820,32'h00000006,32'h00000000,
32'h00100000,32'h00000000,32'h00000000,32'h08000000,32'h02008020,32'h8280a82c,32'h00000009,32'h00000000
};

rcm_mem_bfu_array='{
32'h80000028,32'h0003fa87,32'h00000000,32'h00000000,
32'ha0000028,32'h0003fa97,32'h00000000,32'h00000000,
32'hc0000028,32'h0003faa7,32'h00000000,32'h00000000,
32'he0000028,32'h0003fab7,32'h00000000,32'h00000000,
32'he0000010,32'h0003ffff,32'h00000000,32'h00000000,
32'h0000002a,32'h00016112,32'h00000000,32'h00000000,
32'h4000002a,32'h00016932,32'h00000000,32'h00000000,
32'h8000002a,32'h00017152,32'h00000000,32'h00000000,
32'hc000002a,32'h00017972,32'h00000000,32'h00000000,
32'h00000028,32'h0003f820,32'h00000000,32'h00000000,
32'h00000010,32'h0003fa81,32'h00000000,32'h00000000,
32'h00000010,32'h0003fa91,32'h00000000,32'h00000000,
32'h80000028,32'h0003f860,32'h00000000,32'h00000000,
32'h20000009,32'h0003fc38,32'h00000000,32'h00000000,
32'hd1010404,32'h0003fff9,32'h00000000,32'h00000000,
32'h40000010,32'h0003f839,32'h00000000,32'h00000000,
32'h80000010,32'h0003f829,32'h00000000,32'h00000000,
32'h9101fc24,32'h00022ff0,32'h00000000,32'h00000000,
32'hd0c20004,32'h0003fc70,32'h00000000,32'h00000000,
32'h00000028,32'h0003fae5,32'h00000000,32'h00000000,
32'h20000028,32'h0003faf5,32'h00000000,32'h00000000,
32'h40000028,32'h0003fac5,32'h00000000,32'h00000000,
32'h60000028,32'h0003fad5,32'h00000000,32'h00000000
};

rcm_mem_route_array='{
32'h0fffffff,32'h00000000,32'h00000000,32'h00000000,
32'h00c10100,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd6ac,32'h00000000,32'h00000000,32'h00000000,
32'h00200508,32'h00000000,32'h00000000,32'h00000000
};

rcm_mem_mem_ctrl_array='{
32'h00000001,32'h00000000,32'h1e0001e0,32'h00000000,
32'h00000001,32'h00000000,32'hfe0001e0,32'h00000007,
32'h00000001,32'h00000000,32'h7e0001e0,32'h00000000
};
