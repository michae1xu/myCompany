#define TDES_ECB_DC_TDES_ECB_DC_STR_ADDR 0
#define TDES_ECB_DC_TDES_ECB_DC_END_ADDR 1
#define TDES_ECB_DC_TDES_ECB_DC_CACHE_NUM 12

rcm_mem_rlm_array='{
0xc0200400 0x20040400 0x040400c0 0xffffa000 
0x00001402 0x00000000 0x00000000 0xffff20a0
};

rcm_mem_rcu_array='{
32'h00000000,32'h00050008,32'h00059800,32'h00000000,32'h00000000,32'h00000000,32'h0000fe00,32'h00000000,
32'h00000000,32'h00000000,32'h00008000,32'h00000000,32'h00000000,32'h00000000,32'h0000fe00,32'h00000000,
32'h00000000,32'h00050008,32'h00049800,32'h00000000,32'h00000000,32'h00000000,32'h0000fe00,32'h00000000,
32'h00000041,32'h02040008,32'h00039000,32'h00000000,32'h00000000,32'h00000000,32'h0000fe03,32'h00000000,
32'h00000042,32'h01030008,32'h41028800,32'h00040000,32'h02800000,32'h80401808,32'h0000fe00,32'h00000000,
32'h00200000,32'h00000000,32'h00008000,32'h00000000,32'h00000000,32'h00000000,32'h0000fe00,32'h00000000
};

rcm_mem_bfu_array='{
32'he0000010,32'h0003ffff,32'h00000000,32'h00000000,
32'h00000028,32'h0003fa8c,32'h00000000,32'h00000000,
32'h20000028,32'h0003fa9c,32'h00000000,32'h00000000,
32'h10906004,32'h0003f820,32'h00000000,32'h00000000,
32'h10014004,32'h0003f942,32'h00000000,32'h00000000,
32'h0000002a,32'h000162d4,32'h00000000,32'h00000000,
32'h80000009,32'h0003fad5,32'h00000000,32'h00000000
};

rcm_mem_route_array='{
32'h0fffffff,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd62d,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd021,32'h00000000,32'h00000000,32'h00000000,
32'h0000007f,32'h00000000,32'h00000000,32'h00000000,
32'h0fffc284,32'h00000000,32'h00000000,32'h00000000,
32'h0fffff86,32'h00000000,32'h00000000,32'h00000000,
32'h0fffc488,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd62c,32'h00000000,32'h00000000,32'h00000000,
32'h0fffc080,32'h00000000,32'h00000000,32'h00000000,
32'h0ffff061,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd0a0,32'h00000000,32'h00000000,32'h00000000,
32'h0fffdebc,32'h00000000,32'h00000000,32'h00000000
};

rcm_mem_mem_ctrl_array='{
32'h00000001,32'h00000000,32'h000001e0,32'h00000020,
32'h00000001,32'h00000000,32'h200001e0,32'h00000000,
32'h00000001,32'h00000000,32'h020001e0,32'h00000020
};

