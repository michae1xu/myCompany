
`define des_STR_ADDR 0
`define des_END_ADDR 0
`define des_CACHE_NUM 6
rcm_mem_array='{
32'hc0200400,32'h00140400,32'h00000000,32'hffff6000
};
rcm_mem_rcu_array='{
32'h00000000,32'h00000000,32'h00048000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,
32'h00000000,32'h00010008,32'h00008800,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,
32'h00000041,32'h02040008,32'h00039000,32'h00000000,32'h00000000,32'h00000000,32'h00000003,32'h00000000,
32'h00000002,32'h01030008,32'h41029800,32'h00040000,32'h02800000,32'h80401808,32'h00000000,32'h00000000,
32'h00000000,32'h00000000,32'h0001a000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,
32'h00200000,32'h00000000,32'h00008000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000
};

rcm_mem_bfu_array='{
32'he0000010,32'h0003ffff,32'h00000000,32'h00000000,
32'h00000028,32'h0003fa8c,32'h00000000,32'h00000000,
32'h20000010,32'h0003fa9c,32'h00000000,32'h00000000,
32'h10906004,32'h0003f820,32'h00000000,32'h00000000,
32'h10014004,32'h0003f942,32'h00000000,32'h00000000,
32'h0000002a,32'h00016ac4,32'h00000000,32'h00000000,
32'h80000009,32'h0003fad5,32'h00000000,32'h00000000
};

rcm_mem_route_array='{
32'h0fffffff,32'h00000000,32'h00000000,32'h00000000,
32'h0ffff0e0,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd0a0,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd6ac,32'h00000000,32'h00000000,32'h00000000,
32'h0fffc284,32'h00000000,32'h00000000,32'h00000000,
32'h0fffff86,32'h00000000,32'h00000000,32'h00000000,
32'h0fffc409,32'h00000000,32'h00000000,32'h00000000,
32'h0fffd62c,32'h00000000,32'h00000000,32'h00000000,
32'h0fffc080,32'h00000000,32'h00000000,32'h00000000,
32'h0fffdebc,32'h00000000,32'h00000000,32'h00000000
};

rcm_mem_mem_ctrl_array='{
32'h00000001,32'h00000000,32'h000001e0,32'h00000020,
32'h00000001,32'h00000000,32'h3e0001e0,32'h00000026,
32'h00000001,32'h00000000,32'h020001e0,32'h00000020
};
